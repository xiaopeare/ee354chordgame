module /Users/xiaolei/Desktop/letters/error_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=11'b00000000000) && ({row_reg, col_reg}<11'b00000000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000000110)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00000000111) && ({row_reg, col_reg}<11'b00000011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000011011)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}>=11'b00000011100) && ({row_reg, col_reg}<11'b00000100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000100001)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}>=11'b00000100010) && ({row_reg, col_reg}<11'b00000101001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000101001)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00000101010) && ({row_reg, col_reg}<11'b00000110101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000110101)) color_data = 12'b110110111001;

		if(({row_reg, col_reg}>=11'b00000110110) && ({row_reg, col_reg}<11'b00001000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001000100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00001000101) && ({row_reg, col_reg}<11'b00001100111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001100111)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00001101000) && ({row_reg, col_reg}<11'b00001101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001101111)) color_data = 12'b110110111001;

		if(({row_reg, col_reg}>=11'b00001110000) && ({row_reg, col_reg}<11'b00010000001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010000001)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00010000010) && ({row_reg, col_reg}<11'b00010010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010010110)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00010010111) && ({row_reg, col_reg}<11'b00010011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010011010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b00010011011)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00010011100) && ({row_reg, col_reg}<11'b00010101101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010101101)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00010101110) && ({row_reg, col_reg}<11'b00010110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010110001)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b00010110010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00010110011) && ({row_reg, col_reg}<11'b00010110111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010110111)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b00010111000) && ({row_reg, col_reg}<11'b00011000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011000011)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00011000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b00011000101) && ({row_reg, col_reg}<11'b00011000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00011000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b00011001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b00011001001) && ({row_reg, col_reg}<11'b00011001100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00011001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00011001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00011001110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=11'b00011001111) && ({row_reg, col_reg}<11'b00011011101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011011101)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00011011110) && ({row_reg, col_reg}<11'b00011100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011100011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b00011100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011100101)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00011100110) && ({row_reg, col_reg}<11'b00011101011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011101011)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00011101100) && ({row_reg, col_reg}<11'b00011110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011110000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b00011110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011110010)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}==11'b00011110011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011110100)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b00011110101) && ({row_reg, col_reg}<11'b00100000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100000101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00100000111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00100001000)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b00100001001) && ({row_reg, col_reg}<11'b00100001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100001100)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00100001101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b00100001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00100001111)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b00100010000) && ({row_reg, col_reg}<11'b00100010011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100010011)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100010100) && ({row_reg, col_reg}<11'b00100011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100011010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b00100011011)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}==11'b00100011100)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00100011101) && ({row_reg, col_reg}<11'b00100100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100100000)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100100001) && ({row_reg, col_reg}<11'b00100100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100100011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00100100100) && ({row_reg, col_reg}<11'b00100101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100101110)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100101111) && ({row_reg, col_reg}<11'b00100110010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100110010)) color_data = 12'b110110111010;

		if(({row_reg, col_reg}>=11'b00100110011) && ({row_reg, col_reg}<11'b00101000000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101000000)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00101000001) && ({row_reg, col_reg}<11'b00101000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101000110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00101000111)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==11'b00101001000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101001001)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b00101001010)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00101001011)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00101001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101001101)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00101001110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00101001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101010000)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b00101010001) && ({row_reg, col_reg}<11'b00101011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101011011)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00101011100) && ({row_reg, col_reg}<11'b00101011110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101011110)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b00101011111) && ({row_reg, col_reg}<11'b00101100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101100100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00101100101) && ({row_reg, col_reg}<11'b00101101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101101110)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}>=11'b00101101111) && ({row_reg, col_reg}<11'b00101110011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101110011)) color_data = 12'b110110111010;

		if(({row_reg, col_reg}>=11'b00101110100) && ({row_reg, col_reg}<11'b00110000000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110000000)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}==11'b00110000001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110000010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00110000011) && ({row_reg, col_reg}<11'b00110000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110000111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b00110001000) && ({row_reg, col_reg}<11'b00110001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110001010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00110001011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00110001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110001101)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00110001110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00110001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110010000)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b00110010001) && ({row_reg, col_reg}<11'b00110010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110010011)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b00110010100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00110010101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00110010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b00110011000)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b00110011001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00110011010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00110011011) && ({row_reg, col_reg}<11'b00110011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110011101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00110011110)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b00110011111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00110100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00110100010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b00110100011) && ({row_reg, col_reg}<11'b00110100110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110100110)) color_data = 12'b101110101000;
		if(({row_reg, col_reg}==11'b00110100111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00110101000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00110101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b00110101011)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00110101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110101101)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b00110101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110101111)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00110110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110110001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00110110010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00110110011)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00110110100)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==11'b00110110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b00110110111)) color_data = 12'b101010000111;

		if(({row_reg, col_reg}>=11'b00110111000) && ({row_reg, col_reg}<11'b00111000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111000100)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b00111000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00111000111)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b00111001000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b00111001001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111001010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00111001011)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b00111001100)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b00111001101)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00111001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b00111001111) && ({row_reg, col_reg}<11'b00111010001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111010001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00111010010)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==11'b00111010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00111010100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00111010101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00111010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111010111)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==11'b00111011000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00111011001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00111011010) && ({row_reg, col_reg}<11'b00111011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111011100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00111011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00111011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00111011111)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b00111100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111100001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00111100010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00111100011)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00111100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111100101)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==11'b00111100110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00111100111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00111101000)) color_data = 12'b101110101000;
		if(({row_reg, col_reg}==11'b00111101001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00111101010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00111101011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00111101100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00111101101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b00111101110) && ({row_reg, col_reg}<11'b00111110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111110000)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00111110001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b00111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00111110011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b00111110100)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00111110101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111110110)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==11'b00111110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00111111000)) color_data = 12'b101110011000;

		if(({row_reg, col_reg}>=11'b00111111001) && ({row_reg, col_reg}<11'b01000000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000000011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01000000100) && ({row_reg, col_reg}<11'b01000000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b01000000110) && ({row_reg, col_reg}<11'b01000001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01000001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01000001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01000001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01000001011)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01000001100)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}==11'b01000001101)) color_data = 12'b110010011001;
		if(({row_reg, col_reg}==11'b01000001110)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}>=11'b01000001111) && ({row_reg, col_reg}<11'b01000010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000010010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01000010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01000010100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01000010101) && ({row_reg, col_reg}<11'b01000010111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000010111)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01000011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b01000011001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01000011010) && ({row_reg, col_reg}<11'b01000011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000011100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01000011101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01000011110)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}>=11'b01000011111) && ({row_reg, col_reg}<11'b01000100010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000100010)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01000100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01000100100)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01000100101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01000100110)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==11'b01000100111)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01000101000) && ({row_reg, col_reg}<11'b01000101011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000101011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01000101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01000101101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01000101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000101111)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01000110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000110001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01000110010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01000110011)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01000110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000110101)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01000110110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000110111)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==11'b01000111000)) color_data = 12'b100001100101;

		if(({row_reg, col_reg}>=11'b01000111001) && ({row_reg, col_reg}<11'b01001000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001000101)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==11'b01001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001000111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01001001000)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01001001001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001001010)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01001001011)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01001001100) && ({row_reg, col_reg}<11'b01001010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001010010)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01001010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01001010100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01001010101)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01001010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001010111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01001011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01001011001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01001011010) && ({row_reg, col_reg}<11'b01001011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001011100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01001011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001011110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b01001011111) && ({row_reg, col_reg}<11'b01001100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001100001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01001100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b01001100100)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01001100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01001100110)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01001100111)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01001101000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001101001)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}==11'b01001101010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01001101011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001101100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01001101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b01001101110) && ({row_reg, col_reg}<11'b01001110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001110001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01001110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01001110011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01001110100) && ({row_reg, col_reg}<11'b01001110110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001110110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01001110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001111000)) color_data = 12'b100101110110;

		if(({row_reg, col_reg}>=11'b01001111001) && ({row_reg, col_reg}<11'b01010000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010000011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01010000100) && ({row_reg, col_reg}<11'b01010000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01010000111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01010001000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010001001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01010001010)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==11'b01010001011)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01010001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010001101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01010001110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==11'b01010001111)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01010010000) && ({row_reg, col_reg}<11'b01010010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010010010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01010010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01010010100) && ({row_reg, col_reg}<11'b01010010111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010010111)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01010011000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01010011001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01010011010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01010011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010011100)) color_data = 12'b101010010111;
		if(({row_reg, col_reg}==11'b01010011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010011110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01010011111) && ({row_reg, col_reg}<11'b01010100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010100001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01010100010)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==11'b01010100011)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01010100100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01010100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010100110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b01010100111) && ({row_reg, col_reg}<11'b01010101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010101100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01010101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01010101110) && ({row_reg, col_reg}<11'b01010110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010110001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01010110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01010110011) && ({row_reg, col_reg}<11'b01010110101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010110101)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b01010110110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01010110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01010111000)) color_data = 12'b101110011000;

		if(({row_reg, col_reg}>=11'b01010111001) && ({row_reg, col_reg}<11'b01011000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b01011000011) && ({row_reg, col_reg}<11'b01011000101)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01011000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01011000111)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01011001000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011001001)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b01011001010)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01011001011)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01011001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011001101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01011001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01011001111)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01011010000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011010001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01011010010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01011010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01011010100)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b01011010101) && ({row_reg, col_reg}<11'b01011011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011011100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01011011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01011011110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b01011011111) && ({row_reg, col_reg}<11'b01011100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011100001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01011100010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011100011)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01011100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01011100110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}>=11'b01011100111) && ({row_reg, col_reg}<11'b01011101011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011101011)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01011101100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01011101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01011101110) && ({row_reg, col_reg}<11'b01011110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011110001)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01011110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01011110011) && ({row_reg, col_reg}<11'b01011110111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011110111)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01011111000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011111001)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b01011111010) && ({row_reg, col_reg}<11'b01100000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01100000111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01100001000) && ({row_reg, col_reg}<11'b01100001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100001010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01100001011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100001100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01100001101)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01100001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01100001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100010000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01100010001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100010010)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01100010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01100010100) && ({row_reg, col_reg}<11'b01100010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100010110)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b01100010111) && ({row_reg, col_reg}<11'b01100011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100011010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01100011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100011100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01100011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01100011110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01100011111) && ({row_reg, col_reg}<11'b01100100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01100100110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01100100111)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b01100101000) && ({row_reg, col_reg}<11'b01100101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100101100)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01100101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01100101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100101111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01100110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100110001)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==11'b01100110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01100110011) && ({row_reg, col_reg}<11'b01100110101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b01100110101) && ({row_reg, col_reg}<11'b01100110111)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b01100110111) && ({row_reg, col_reg}<11'b01101000010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101000010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01101000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101000100)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01101000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01101000111)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}>=11'b01101001000) && ({row_reg, col_reg}<11'b01101001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101001010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01101001011) && ({row_reg, col_reg}<11'b01101001101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101001101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01101001110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01101001111)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01101010000) && ({row_reg, col_reg}<11'b01101010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101010010)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01101010100) && ({row_reg, col_reg}<11'b01101011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101011100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01101011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101011110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01101011111) && ({row_reg, col_reg}<11'b01101100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101100011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01101100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101100101)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01101100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01101100111)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01101101000) && ({row_reg, col_reg}<11'b01101101010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101101010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01101101011)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==11'b01101101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101101101)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01101101110)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01101101111)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}==11'b01101110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101110001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01101110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01101110011) && ({row_reg, col_reg}<11'b01101110110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101110110)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b01101110111) && ({row_reg, col_reg}<11'b01110000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110000100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01110000101)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01110001000)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01110001001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01110001010)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01110001011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01110001100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01110001101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b01110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110001111)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}>=11'b01110010000) && ({row_reg, col_reg}<11'b01110010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110010010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01110010011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01110010100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01110010101) && ({row_reg, col_reg}<11'b01110010111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110010111)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}>=11'b01110011000) && ({row_reg, col_reg}<11'b01110011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110011010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01110011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110011100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01110011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110011110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01110011111)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01110100000) && ({row_reg, col_reg}<11'b01110100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110100100)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b01110100101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01110100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01110100111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01110101000)) color_data = 12'b101110101000;
		if(({row_reg, col_reg}==11'b01110101001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110101010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01110101011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01110101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=11'b01110101101) && ({row_reg, col_reg}<11'b01110101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110101111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01110110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110110001)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==11'b01110110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110110011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01110110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110110101)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b01110110110) && ({row_reg, col_reg}<11'b01111000001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111000001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01111000010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111000011)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01111000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01111000110) && ({row_reg, col_reg}<11'b01111001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=11'b01111001001) && ({row_reg, col_reg}<11'b01111001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111001011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=11'b01111001100) && ({row_reg, col_reg}<11'b01111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111010000)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01111010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01111010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111010101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=11'b01111010110) && ({row_reg, col_reg}<11'b01111011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111011010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01111011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01111011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111011101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01111011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01111100000)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01111100001) && ({row_reg, col_reg}<11'b01111100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111100011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01111100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111100101)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01111100110)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==11'b01111100111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01111101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111101010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01111101011)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01111101100)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01111101101) && ({row_reg, col_reg}<11'b01111101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111101111)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==11'b01111110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01111110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111110010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==11'b01111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111110100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=11'b01111110101) && ({row_reg, col_reg}<11'b01111111010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111111010)) color_data = 12'b110110101001;





		if(({row_reg, col_reg}>=11'b01111111011) && ({row_reg, col_reg}<=11'b10011111011)) color_data = 12'b110010101001;
	end
endmodule