module /Users/xiaolei/Desktop/letters/lvl2_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=11'b00000000000) && ({row_reg, col_reg}<11'b00000000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000000110)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00000000111) && ({row_reg, col_reg}<11'b00000001011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000001011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00000001100) && ({row_reg, col_reg}<11'b00000011101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000011101)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00000011110) && ({row_reg, col_reg}<11'b00000100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000100001)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00000100010) && ({row_reg, col_reg}<11'b00000101000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000101000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00000101001) && ({row_reg, col_reg}<11'b00000110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000110001)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b00000110010) && ({row_reg, col_reg}<11'b00001000000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001000000)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b00001000001) && ({row_reg, col_reg}<11'b00001001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001001010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00001001011) && ({row_reg, col_reg}<11'b00001010100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001010100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00001010101) && ({row_reg, col_reg}<11'b00001011000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001011000)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b00001011001) && ({row_reg, col_reg}<11'b00001011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001011011)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00001011100) && ({row_reg, col_reg}<11'b00001100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001100100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b00001100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001100110)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00001100111) && ({row_reg, col_reg}<11'b00001101101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001101101)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00001101110) && ({row_reg, col_reg}<11'b00001110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001110000)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b00001110001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00001110010) && ({row_reg, col_reg}<11'b00001110101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001110101)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b00001110110) && ({row_reg, col_reg}<11'b00001111010)) color_data = 12'b110010101001;

		if(({row_reg, col_reg}>=11'b00001111010) && ({row_reg, col_reg}<11'b00010000000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00010000000) && ({row_reg, col_reg}<11'b00010000010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010000010)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}==11'b00010000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b00010000100) && ({row_reg, col_reg}<11'b00010000110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00010000110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00010000111) && ({row_reg, col_reg}<11'b00010001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010001100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b00010001101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010001110)) color_data = 12'b101110101000;
		if(({row_reg, col_reg}>=11'b00010001111) && ({row_reg, col_reg}<11'b00010010001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b00010010001) && ({row_reg, col_reg}<11'b00010011000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b00010011000) && ({row_reg, col_reg}<11'b00010011010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00010011010)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b00010011011) && ({row_reg, col_reg}<11'b00010011101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010011101)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b00010011110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010011111)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00010100000) && ({row_reg, col_reg}<11'b00010100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010100101)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}==11'b00010100110)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00010100111) && ({row_reg, col_reg}<11'b00010110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010110001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00010110010)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b00010110011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00010110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00010110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b00010110110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00010110111)) color_data = 12'b101110011000;

		if(({row_reg, col_reg}>=11'b00010111000) && ({row_reg, col_reg}<11'b00011000010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011000010)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00011000011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00011000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b00011000101) && ({row_reg, col_reg}<11'b00011000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00011000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b00011001000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00011001001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00011001010) && ({row_reg, col_reg}<11'b00011001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011001100)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==11'b00011001101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00011001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b00011001111) && ({row_reg, col_reg}<11'b00011010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b00011010001) && ({row_reg, col_reg}<11'b00011010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00011010011)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b00011010100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011010101)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00011010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b00011010111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00011011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00011011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00011011010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00011011011)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00011011100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00011011101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00011011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00011011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00011100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00011100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b00011100010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00011100011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00011100100)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00011100101) && ({row_reg, col_reg}<11'b00011110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011110000)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00011110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00011110010)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00011110011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00011110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011110101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00011110110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00011110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00011111000)) color_data = 12'b101010011000;

		if(({row_reg, col_reg}>=11'b00011111001) && ({row_reg, col_reg}<11'b00100000000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100000000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00100000001) && ({row_reg, col_reg}<11'b00100000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100000100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00100000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00100000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=11'b00100000111) && ({row_reg, col_reg}<11'b00100001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100001110)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==11'b00100001111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00100010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00100010001)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==11'b00100010010)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b00100010011) && ({row_reg, col_reg}<11'b00100010111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100010111)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00100011000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00100011001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b00100011010) && ({row_reg, col_reg}<11'b00100011110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100011110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00100011111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00100100000)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=11'b00100100001) && ({row_reg, col_reg}<11'b00100100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100100011)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==11'b00100100100)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}>=11'b00100100101) && ({row_reg, col_reg}<11'b00100101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100101111)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00100110000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00100110001)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00100110010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100110011) && ({row_reg, col_reg}<11'b00100110111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100110111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00100111000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00100111001)) color_data = 12'b101110011001;

		if(({row_reg, col_reg}>=11'b00100111010) && ({row_reg, col_reg}<11'b00101000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101000100)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==11'b00101000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00101000110)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b00101000111) && ({row_reg, col_reg}<11'b00101001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101001010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00101001011) && ({row_reg, col_reg}<11'b00101001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101001111)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00101010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00101010001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00101010010)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b00101010011) && ({row_reg, col_reg}<11'b00101010111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101010111)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==11'b00101011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00101011001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00101011010) && ({row_reg, col_reg}<11'b00101011110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101011110)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b00101011111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00101100000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b00101100001) && ({row_reg, col_reg}<11'b00101100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101100100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00101100101) && ({row_reg, col_reg}<11'b00101101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101101111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00101110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00101110001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00101110010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101110011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00101110100) && ({row_reg, col_reg}<11'b00101110111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101110111)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00101111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00101111001)) color_data = 12'b101110011000;

		if(({row_reg, col_reg}>=11'b00101111010) && ({row_reg, col_reg}<11'b00110000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00110000110)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}>=11'b00110000111) && ({row_reg, col_reg}<11'b00110001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110001111)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b00110010000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00110010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110010010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00110010011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00110010100) && ({row_reg, col_reg}<11'b00110010111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110010111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00110011000)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==11'b00110011001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110011010)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==11'b00110011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110011100)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00110011101) && ({row_reg, col_reg}<11'b00110011111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110100000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b00110100001) && ({row_reg, col_reg}<11'b00110100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110100100)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00110100101) && ({row_reg, col_reg}<11'b00110101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110101111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b00110110000) && ({row_reg, col_reg}<11'b00110110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b00110110010) && ({row_reg, col_reg}<11'b00110110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110110100)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00110110101) && ({row_reg, col_reg}<11'b00110110111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110110111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00110111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110111001)) color_data = 12'b101110101001;

		if(({row_reg, col_reg}>=11'b00110111010) && ({row_reg, col_reg}<11'b00111000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00111000110)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b00111000111) && ({row_reg, col_reg}<11'b00111001011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111001011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00111001100) && ({row_reg, col_reg}<11'b00111010000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111010000)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00111010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00111010010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00111010011) && ({row_reg, col_reg}<11'b00111010111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b00111011000)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00111011001)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b00111011010) && ({row_reg, col_reg}<11'b00111011110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111011110)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b00111011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00111100000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b00111100001) && ({row_reg, col_reg}<11'b00111100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111100101)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00111100110) && ({row_reg, col_reg}<11'b00111101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111101110)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b00111101111)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}==11'b00111110000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00111110001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b00111110010) && ({row_reg, col_reg}<11'b00111110110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111110110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00111110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00111111000)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=11'b00111111001) && ({row_reg, col_reg}<11'b00111111011)) color_data = 12'b110010101001;

		if(({row_reg, col_reg}==11'b00111111011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01000000000) && ({row_reg, col_reg}<11'b01000000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01000000110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01000000111) && ({row_reg, col_reg}<11'b01000001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000001010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01000001011) && ({row_reg, col_reg}<11'b01000001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000001111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01000010000)) color_data = 12'b110010011001;
		if(({row_reg, col_reg}==11'b01000010001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==11'b01000010010)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=11'b01000010011) && ({row_reg, col_reg}<11'b01000010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000010110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01000010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01000011000)) color_data = 12'b110010011001;
		if(({row_reg, col_reg}>=11'b01000011001) && ({row_reg, col_reg}<11'b01000011111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01000100000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01000100001) && ({row_reg, col_reg}<11'b01000100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000100011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01000100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000100101)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01000100110) && ({row_reg, col_reg}<11'b01000110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000110100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01000110101)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=11'b01000110110) && ({row_reg, col_reg}<11'b01000111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01000111000)) color_data = 12'b101010000111;

		if(({row_reg, col_reg}>=11'b01000111001) && ({row_reg, col_reg}<11'b01001000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001000110)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}>=11'b01001000111) && ({row_reg, col_reg}<11'b01001001011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001001011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01001001100) && ({row_reg, col_reg}<11'b01001001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001001110)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b01001001111) && ({row_reg, col_reg}<11'b01001010001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001010001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01001010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001010011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01001010100) && ({row_reg, col_reg}<11'b01001010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001010110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01001010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=11'b01001011000) && ({row_reg, col_reg}<11'b01001011111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001100000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01001100001)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b01001100010) && ({row_reg, col_reg}<11'b01001100111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001100111)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b01001101000) && ({row_reg, col_reg}<11'b01001101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001101111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01001110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001110001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01001110010)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b01001110011) && ({row_reg, col_reg}<11'b01001110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001110110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01001110111)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01001111000)) color_data = 12'b110010101010;

		if(({row_reg, col_reg}>=11'b01001111001) && ({row_reg, col_reg}<11'b01010000000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010000000)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b01010000001) && ({row_reg, col_reg}<11'b01010000011)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b01010000011) && ({row_reg, col_reg}<11'b01010000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010000110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01010000111) && ({row_reg, col_reg}<11'b01010001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010001010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01010001011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010001100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01010001101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==11'b01010001110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01010001111) && ({row_reg, col_reg}<11'b01010010001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010010001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01010010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01010010011)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=11'b01010010100) && ({row_reg, col_reg}<11'b01010010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010010111)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01010011000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010011001)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b01010011010) && ({row_reg, col_reg}<11'b01010011111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01010100000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01010100001) && ({row_reg, col_reg}<11'b01010100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010100011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01010100100) && ({row_reg, col_reg}<11'b01010100110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010100110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01010100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01010101000)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}>=11'b01010101001) && ({row_reg, col_reg}<11'b01010101101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010101101)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}>=11'b01010101110) && ({row_reg, col_reg}<11'b01010110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010110000)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01010110001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01010110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01010110011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b01010110100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01010110101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01010110110) && ({row_reg, col_reg}<11'b01010111011)) color_data = 12'b110010101001;

		if(({row_reg, col_reg}==11'b01010111011)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b01011000000) && ({row_reg, col_reg}<11'b01011000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011000011)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01011000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b01011000110)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b01011000111) && ({row_reg, col_reg}<11'b01011001001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01011001001) && ({row_reg, col_reg}<11'b01011001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011001100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01011001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01011001110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01011001111) && ({row_reg, col_reg}<11'b01011010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01011010011)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==11'b01011010100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011010101)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01011010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01011010111) && ({row_reg, col_reg}<11'b01011011111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011011111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01011100000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b01011100001) && ({row_reg, col_reg}<11'b01011100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011100100)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01011100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011100110)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01011100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01011101000)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}>=11'b01011101001) && ({row_reg, col_reg}<11'b01011101011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011101011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01011101100) && ({row_reg, col_reg}<11'b01011101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011101111)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01011110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01011110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01011110010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01011110011) && ({row_reg, col_reg}<11'b01011110111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011110111)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==11'b01011111000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01011111001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01011111010)) color_data = 12'b110010111010;

		if(({row_reg, col_reg}==11'b01011111011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100000000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01100000001) && ({row_reg, col_reg}<11'b01100000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01100000110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01100000111) && ({row_reg, col_reg}<11'b01100001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100001010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01100001011)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01100001100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01100001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01100001110) && ({row_reg, col_reg}<11'b01100010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100010010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01100010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01100010100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100010101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01100010110)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01100010111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100011000)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01100011001) && ({row_reg, col_reg}<11'b01100011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100011011)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b01100011100) && ({row_reg, col_reg}<11'b01100011111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01100100000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01100100001)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b01100100010) && ({row_reg, col_reg}<11'b01100100110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100100110)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01100100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01100101000) && ({row_reg, col_reg}<11'b01100101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100101110)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01100101111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01100110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01100110001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01100110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01100110011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01100110100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01100110101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100110110)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01100110111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01100111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01100111001)) color_data = 12'b011101010100;

		if(({row_reg, col_reg}>=11'b01100111010) && ({row_reg, col_reg}<11'b01101000000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101000000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01101000001) && ({row_reg, col_reg}<11'b01101000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101000110)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01101000111)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}>=11'b01101001000) && ({row_reg, col_reg}<11'b01101001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101001100)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==11'b01101001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01101001110) && ({row_reg, col_reg}<11'b01101010001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101010001)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01101010010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101010100)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==11'b01101010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01101010110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b01101010111) && ({row_reg, col_reg}<11'b01101011101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101011101)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01101011110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01101100000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b01101100001) && ({row_reg, col_reg}<11'b01101100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101100101)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01101100110)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01101100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01101101000) && ({row_reg, col_reg}<11'b01101101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01101110000)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}>=11'b01101110001) && ({row_reg, col_reg}<11'b01101110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01101110100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01101110101)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01101110110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01101110111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101111000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01101111001)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01101111010)) color_data = 12'b110010101001;

		if(({row_reg, col_reg}==11'b01101111011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01110000000) && ({row_reg, col_reg}<11'b01110000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110000100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01110000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=11'b01110000111) && ({row_reg, col_reg}<11'b01110001001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110001001)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b01110001010) && ({row_reg, col_reg}<11'b01110001100)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01110001100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01110001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110001110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01110001111)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01110010000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01110010001) && ({row_reg, col_reg}<11'b01110010011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110010011)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==11'b01110010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01110010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01110010110)) color_data = 12'b110010011001;
		if(({row_reg, col_reg}==11'b01110010111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110011000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01110011001) && ({row_reg, col_reg}<11'b01110011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110011100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01110011101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110011110)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01110011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110100000)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01110100001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01110100010)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b01110100011) && ({row_reg, col_reg}<11'b01110100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110100101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01110100110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01110100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01110101000) && ({row_reg, col_reg}<11'b01110101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01110110000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=11'b01110110001) && ({row_reg, col_reg}<11'b01110110011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01110110011)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01110110100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01110110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01110110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01110110111) && ({row_reg, col_reg}<11'b01110111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110111001)) color_data = 12'b101010000111;

		if(({row_reg, col_reg}>=11'b01110111010) && ({row_reg, col_reg}<11'b01111000001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111000001)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==11'b01111000010)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01111000011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b01111000100) && ({row_reg, col_reg}<11'b01111000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01111001000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01111001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01111001011) && ({row_reg, col_reg}<11'b01111001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=11'b01111001110) && ({row_reg, col_reg}<11'b01111010000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111010000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01111010001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01111010010)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01111010011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01111010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111010101)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01111010110) && ({row_reg, col_reg}<11'b01111011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111011100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b01111011101) && ({row_reg, col_reg}<11'b01111011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=11'b01111011111) && ({row_reg, col_reg}<11'b01111100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01111100011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01111100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01111100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01111100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=11'b01111101000) && ({row_reg, col_reg}<11'b01111101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111101110)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==11'b01111101111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01111110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111110001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01111110010) && ({row_reg, col_reg}<11'b01111110101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111110101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01111110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b01111110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111111000)) color_data = 12'b100101110110;





		if(({row_reg, col_reg}>=11'b01111111001) && ({row_reg, col_reg}<=11'b10011111011)) color_data = 12'b110010101001;
	end
endmodule