module /Users/xiaolei/Desktop/letters/aug_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=11'b00000000000) && ({row_reg, col_reg}<11'b00000001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000001110)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00000001111) && ({row_reg, col_reg}<11'b00000100010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000100010)) color_data = 12'b110010111001;

		if(({row_reg, col_reg}>=11'b00000100011) && ({row_reg, col_reg}<11'b00001010000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001010000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00001010001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00001010010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00001010011) && ({row_reg, col_reg}<11'b00001010101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001010101)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00001010110) && ({row_reg, col_reg}<11'b00001011001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001011001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00001011010) && ({row_reg, col_reg}<11'b00001011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b00001011100) && ({row_reg, col_reg}<11'b00001011110)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b00001011110) && ({row_reg, col_reg}<11'b00010001001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010001001)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00010001010) && ({row_reg, col_reg}<11'b00010001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010001111)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==11'b00010010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00010010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b00010010010)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}>=11'b00010010011) && ({row_reg, col_reg}<11'b00010011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010011100)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}>=11'b00010011101) && ({row_reg, col_reg}<11'b00010100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010100001)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b00010100010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b00010100011) && ({row_reg, col_reg}<11'b00010100101)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00010100101) && ({row_reg, col_reg}<11'b00010101000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010101000)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b00010101001) && ({row_reg, col_reg}<11'b00011001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011001111)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00011010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00011010001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00011010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b00011010011) && ({row_reg, col_reg}<11'b00011010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011010110)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00011010111) && ({row_reg, col_reg}<11'b00011011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011011100)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b00011011101) && ({row_reg, col_reg}<11'b00011011111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011011111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00011100000) && ({row_reg, col_reg}<11'b00011100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011100011)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}==11'b00011100100)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00011100101) && ({row_reg, col_reg}<11'b00011101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011101100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00011101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00011101110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00011101111)) color_data = 12'b100110000111;

		if(({row_reg, col_reg}>=11'b00011110000) && ({row_reg, col_reg}<11'b00100001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100001110)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b00100001111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00100010000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00100010001)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00100010010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b00100010011)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b00100010100) && ({row_reg, col_reg}<11'b00100010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100010110)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b00100010111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100011000)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100011001) && ({row_reg, col_reg}<11'b00100011101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100011101)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100011110) && ({row_reg, col_reg}<11'b00100101011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100101011)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==11'b00100101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00100101101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00100101110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00100101111)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}>=11'b00100110000) && ({row_reg, col_reg}<11'b00101001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101001010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00101001011) && ({row_reg, col_reg}<11'b00101001101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101001101)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b00101001110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00101001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00101010000)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00101010001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101010010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00101010011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=11'b00101010100) && ({row_reg, col_reg}<11'b00101011000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101011000)) color_data = 12'b101110101000;
		if(({row_reg, col_reg}==11'b00101011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00101011010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==11'b00101011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b00101011100) && ({row_reg, col_reg}<11'b00101011110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00101011110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101011111)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}==11'b00101100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b00101100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00101100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=11'b00101100011) && ({row_reg, col_reg}<11'b00101101000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101101000)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00101101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b00101101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b00101101011) && ({row_reg, col_reg}<11'b00101101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00101101101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00101101110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00101101111)) color_data = 12'b011001010011;

		if(({row_reg, col_reg}>=11'b00101110000) && ({row_reg, col_reg}<11'b00110001101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110001101)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b00110001110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00110001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110010000)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00110010001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b00110010010)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==11'b00110010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b00110010100) && ({row_reg, col_reg}<11'b00110011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110011010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00110011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110011100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00110011101)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b00110011110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110011111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b00110100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110100001)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==11'b00110100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b00110100011) && ({row_reg, col_reg}<11'b00110100111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110100111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00110101000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110101001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00110101010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00110101011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00110101100)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00110101101)) color_data = 12'b010100110010;

		if(({row_reg, col_reg}>=11'b00110101110) && ({row_reg, col_reg}<11'b00111001011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111001011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00111001100) && ({row_reg, col_reg}<11'b00111001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111001110)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==11'b00111001111)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}>=11'b00111010000) && ({row_reg, col_reg}<11'b00111010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111010010)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b00111010011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00111010100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b00111010101) && ({row_reg, col_reg}<11'b00111011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111011010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00111011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00111011100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00111011101) && ({row_reg, col_reg}<11'b00111100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111100001)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00111100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b00111100011) && ({row_reg, col_reg}<11'b00111100111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b00111101000)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}>=11'b00111101001) && ({row_reg, col_reg}<11'b00111101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111101100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00111101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b00111101110)) color_data = 12'b101110011000;

		if(({row_reg, col_reg}>=11'b00111101111) && ({row_reg, col_reg}<11'b01000001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000001100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01000001101)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01000001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01000001111)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b01000010000) && ({row_reg, col_reg}<11'b01000010011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01000010100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01000010101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b01000010110) && ({row_reg, col_reg}<11'b01000011000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01000011000) && ({row_reg, col_reg}<11'b01000011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000011010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01000011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01000011100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=11'b01000011101) && ({row_reg, col_reg}<11'b01000100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000100000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01000100001)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01000100010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=11'b01000100011) && ({row_reg, col_reg}<11'b01000100111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01000101000)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01000101001) && ({row_reg, col_reg}<11'b01000101011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000101011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01000101100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01000101101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01000101110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01000101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000110000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01000110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000110010)) color_data = 12'b110110111001;

		if(({row_reg, col_reg}>=11'b01000110011) && ({row_reg, col_reg}<11'b01001001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001001010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01001001011) && ({row_reg, col_reg}<11'b01001001101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001001101)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01001001110) && ({row_reg, col_reg}<11'b01001010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01001010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b01001010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01001010101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01001010110) && ({row_reg, col_reg}<11'b01001011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001011010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01001011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01001011100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01001011101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001011110)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01001011111) && ({row_reg, col_reg}<11'b01001100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001100001)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01001100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001100011)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b01001100100) && ({row_reg, col_reg}<11'b01001100110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001100110)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01001100111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b01001101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01001101001)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01001101010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001101011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01001101100)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01001101101)) color_data = 12'b011001010100;

		if(({row_reg, col_reg}>=11'b01001101110) && ({row_reg, col_reg}<11'b01010001000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010001000)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01010001001) && ({row_reg, col_reg}<11'b01010001101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==11'b01010001110)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01010001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010010000)) color_data = 12'b110010011001;
		if(({row_reg, col_reg}==11'b01010010001)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}==11'b01010010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010010011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01010010100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01010010101)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01010010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010010111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01010011000) && ({row_reg, col_reg}<11'b01010011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010011010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01010011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010011100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01010011101)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01010011110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01010011111) && ({row_reg, col_reg}<11'b01010100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010100001)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01010100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01010100011) && ({row_reg, col_reg}<11'b01010100110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010100110)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01010100111)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==11'b01010101000)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==11'b01010101001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01010101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01010101011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01010101100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01010101101)) color_data = 12'b110010111001;

		if(({row_reg, col_reg}>=11'b01010101110) && ({row_reg, col_reg}<11'b01011001001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011001001)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01011001010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01011001011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011001100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01011001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01011001110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b01011001111) && ({row_reg, col_reg}<11'b01011010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011010010)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01011010011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01011010101)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=11'b01011010110) && ({row_reg, col_reg}<11'b01011011001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011011001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01011011010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01011011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01011011100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b01011011101) && ({row_reg, col_reg}<11'b01011011111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011011111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01011100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011100001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01011100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01011100011) && ({row_reg, col_reg}<11'b01011100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011100101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01011100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01011100111)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01011101000)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b01011101001) && ({row_reg, col_reg}<11'b01011101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011101111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01011110000) && ({row_reg, col_reg}<11'b01011110010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011110010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01011110011)) color_data = 12'b110110111001;

		if(({row_reg, col_reg}>=11'b01011110100) && ({row_reg, col_reg}<11'b01100001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100001100)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01100001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=11'b01100001110) && ({row_reg, col_reg}<11'b01100010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100010010)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01100010011)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01100010100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01100010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01100010110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01100010111) && ({row_reg, col_reg}<11'b01100011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100011011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01100011100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01100011101) && ({row_reg, col_reg}<11'b01100011111)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01100011111) && ({row_reg, col_reg}<11'b01100100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100100001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01100100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01100100011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01100100100) && ({row_reg, col_reg}<11'b01100100110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01100100111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01100101000)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01100101001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01100101010) && ({row_reg, col_reg}<11'b01100101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100101100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01100101101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100101110)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}>=11'b01100101111) && ({row_reg, col_reg}<11'b01100110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100110001)) color_data = 12'b110110111001;

		if(({row_reg, col_reg}>=11'b01100110010) && ({row_reg, col_reg}<11'b01101001001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101001001)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01101001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101001011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01101001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101001101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=11'b01101001110) && ({row_reg, col_reg}<11'b01101010001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101010001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01101010010)) color_data = 12'b110010011001;
		if(({row_reg, col_reg}==11'b01101010011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101010100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01101010101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01101010110)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b01101010111) && ({row_reg, col_reg}<11'b01101011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101011011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01101011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01101011101)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b01101011110) && ({row_reg, col_reg}<11'b01101100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101100000)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01101100001) && ({row_reg, col_reg}<11'b01101100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101100011)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=11'b01101100100) && ({row_reg, col_reg}<11'b01101100110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101100110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01101100111)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==11'b01101101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01101101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01101101010) && ({row_reg, col_reg}<11'b01101101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01101101100)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01101101101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01101101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101101111)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01101110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101110001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01101110010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01101110011)) color_data = 12'b100001100101;

		if(({row_reg, col_reg}>=11'b01101110100) && ({row_reg, col_reg}<11'b01110001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110001010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01110001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01110001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01110001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01110010000)) color_data = 12'b101010010111;
		if(({row_reg, col_reg}==11'b01110010001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110010010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=11'b01110010011) && ({row_reg, col_reg}<11'b01110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=11'b01110010110) && ({row_reg, col_reg}<11'b01110011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110011000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01110011001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01110011010) && ({row_reg, col_reg}<11'b01110011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110011100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01110011101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01110011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01110011111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01110100000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01110100001)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01110100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110100011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01110100100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01110100101)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}==11'b01110100110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01110100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01110101000)) color_data = 12'b101010010111;
		if(({row_reg, col_reg}==11'b01110101001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01110101010) && ({row_reg, col_reg}<11'b01110101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110101100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=11'b01110101101) && ({row_reg, col_reg}<11'b01110101111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=11'b01110101111) && ({row_reg, col_reg}<11'b01110110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110110001)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01110110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01110110011)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b01110110100) && ({row_reg, col_reg}<11'b01110110111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110110111)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b01110111000) && ({row_reg, col_reg}<11'b01111001011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111001011)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01111001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111001101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01111001110)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b01111001111) && ({row_reg, col_reg}<11'b01111010101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111010101)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b01111010110) && ({row_reg, col_reg}<11'b01111011110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111011110)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b01111011111) && ({row_reg, col_reg}<11'b01111100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111100001)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b01111100010) && ({row_reg, col_reg}<11'b01111100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111100101)) color_data = 12'b101010010111;
		if(({row_reg, col_reg}==11'b01111100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01111100111)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=11'b01111101000) && ({row_reg, col_reg}<11'b01111101101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111101101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01111101110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01111101111)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==11'b01111110000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111110001)) color_data = 12'b110010111001;

		if(({row_reg, col_reg}>=11'b01111110010) && ({row_reg, col_reg}<11'b10000100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10000100101)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b10000100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b10000100111)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b10000101000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10000101001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b10000101010) && ({row_reg, col_reg}<11'b10000101101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10000101101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b10000101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b10000101111)) color_data = 12'b101010000111;

		if(({row_reg, col_reg}>=11'b10000110000) && ({row_reg, col_reg}<11'b10001100110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10001100110)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b10001100111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b10001101000)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b10001101001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b10001101010) && ({row_reg, col_reg}<11'b10001101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10001101100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b10001101101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b10001101110)) color_data = 12'b011101010100;

		if(({row_reg, col_reg}>=11'b10001101111) && ({row_reg, col_reg}<11'b10010100010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10010100010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b10010100011) && ({row_reg, col_reg}<11'b10010100110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10010100110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b10010100111)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==11'b10010101000)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b10010101001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b10010101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b10010101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b10010101100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b10010101101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b10010101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10010101111)) color_data = 12'b110010111001;

		if(({row_reg, col_reg}>=11'b10010110000) && ({row_reg, col_reg}<11'b10011100100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10011100100)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b10011100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10011100110)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b10011100111) && ({row_reg, col_reg}<11'b10011101101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b10011101101)) color_data = 12'b110110111010;

		if(({row_reg, col_reg}>=11'b10011101110) && ({row_reg, col_reg}<=11'b10011111011)) color_data = 12'b110010101001;
	end
endmodule