module /Users/xiaolei/Desktop/letters/minor_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}==11'b00000000000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00000000001) && ({row_reg, col_reg}<11'b00000100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00000100011)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}==11'b00000100100)) color_data = 12'b110010111001;

		if(({row_reg, col_reg}>=11'b00000100101) && ({row_reg, col_reg}<11'b00001000101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001000101)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b00001000110) && ({row_reg, col_reg}<11'b00001001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001001110)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00001001111) && ({row_reg, col_reg}<11'b00001010010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001010010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00001010011) && ({row_reg, col_reg}<11'b00001010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001010110)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}>=11'b00001010111) && ({row_reg, col_reg}<11'b00001011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001011010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00001011011) && ({row_reg, col_reg}<11'b00001100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001100011)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b00001100100) && ({row_reg, col_reg}<11'b00001100111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001100111)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00001101000) && ({row_reg, col_reg}<11'b00001110101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00001110101)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b00001110110) && ({row_reg, col_reg}<11'b00010000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b00010000011) && ({row_reg, col_reg}<11'b00010000101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00010000101) && ({row_reg, col_reg}<11'b00010010000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010010000)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00010010001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b00010010010) && ({row_reg, col_reg}<11'b00010010101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010010101)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00010010110) && ({row_reg, col_reg}<11'b00010011111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010011111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00010100000) && ({row_reg, col_reg}<11'b00010100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010100101)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00010100110) && ({row_reg, col_reg}<11'b00010110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010110100)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00010110101) && ({row_reg, col_reg}<11'b00010111010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00010111010)) color_data = 12'b110110111010;

		if(({row_reg, col_reg}>=11'b00010111011) && ({row_reg, col_reg}<11'b00011000001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011000001)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b00011000010) && ({row_reg, col_reg}<11'b00011000100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00011000100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00011000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00011000110)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=11'b00011000111) && ({row_reg, col_reg}<11'b00011001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011001010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00011001011) && ({row_reg, col_reg}<11'b00011001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011001110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=11'b00011001111) && ({row_reg, col_reg}<11'b00011010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00011010001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==11'b00011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b00011010011)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=11'b00011010100) && ({row_reg, col_reg}<11'b00011010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b00011010110) && ({row_reg, col_reg}<11'b00011011000)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=11'b00011011000) && ({row_reg, col_reg}<11'b00011011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011011010)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00011011011) && ({row_reg, col_reg}<11'b00011100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011100000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b00011100001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00011100010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00011100011) && ({row_reg, col_reg}<11'b00011101001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b00011101001) && ({row_reg, col_reg}<11'b00011101011)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b00011101011) && ({row_reg, col_reg}<11'b00100000000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100000000)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100000001) && ({row_reg, col_reg}<11'b00100000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100000011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00100000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00100000101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00100000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00100000111)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}>=11'b00100001000) && ({row_reg, col_reg}<11'b00100001011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100001011)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b00100001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100001101)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00100001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00100001111)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b00100010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00100010001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00100010010)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b00100010011) && ({row_reg, col_reg}<11'b00100010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100010110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00100010111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=11'b00100011000) && ({row_reg, col_reg}<11'b00100011101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100011101)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100011110) && ({row_reg, col_reg}<11'b00100101011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100101011)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100101100) && ({row_reg, col_reg}<11'b00100101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100101110)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100101111) && ({row_reg, col_reg}<11'b00100110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100110001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100110010) && ({row_reg, col_reg}<11'b00100110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100110100)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}==11'b00100110101)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00100110110) && ({row_reg, col_reg}<11'b00100111000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00100111000)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==11'b00100111001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b00100111010)) color_data = 12'b110010101001;

		if(({row_reg, col_reg}==11'b00100111011)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b00101000000) && ({row_reg, col_reg}<11'b00101000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00101000101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00101000110)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==11'b00101000111)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}>=11'b00101001000) && ({row_reg, col_reg}<11'b00101001101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101001101)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b00101001110)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00101001111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00101010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00101010001)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b00101010010) && ({row_reg, col_reg}<11'b00101010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}>=11'b00101010110) && ({row_reg, col_reg}<11'b00101011000)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b00101011000) && ({row_reg, col_reg}<11'b00101011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101011011)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b00101011100) && ({row_reg, col_reg}<11'b00101011111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101011111)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b00101100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101100001)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b00101100010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101100011)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b00101100100) && ({row_reg, col_reg}<11'b00101101001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101101001)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b00101101010) && ({row_reg, col_reg}<11'b00101101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101101100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b00101101101) && ({row_reg, col_reg}<11'b00101110111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101110111)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b00101111000) && ({row_reg, col_reg}<11'b00101111010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00101111010)) color_data = 12'b110010111010;

		if(({row_reg, col_reg}>=11'b00101111011) && ({row_reg, col_reg}<11'b00110000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110000101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00110000110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b00110001000) && ({row_reg, col_reg}<11'b00110001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110001010)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}>=11'b00110001011) && ({row_reg, col_reg}<11'b00110001101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110001110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00110001111)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==11'b00110010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b00110010001) && ({row_reg, col_reg}<11'b00110010100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110010100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00110010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110010110)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==11'b00110010111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=11'b00110011000) && ({row_reg, col_reg}<11'b00110011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110011010)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00110011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b00110011101)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b00110011110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00110011111)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b00110100000) && ({row_reg, col_reg}<11'b00110100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110100010)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b00110100011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00110100100) && ({row_reg, col_reg}<11'b00110100110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110100110)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b00110100111) && ({row_reg, col_reg}<11'b00110101001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110101001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00110101010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00110101011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00110101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110101101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00110101110)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00110101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110110000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b00110110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00110110010)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00110110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b00110110101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b00110110110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00110110111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00110111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00110111001)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00110111010)) color_data = 12'b101010000111;

		if(({row_reg, col_reg}==11'b00110111011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111000000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b00111000001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111000010)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==11'b00111000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00111000101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b00111000110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00111000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00111001000)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=11'b00111001001) && ({row_reg, col_reg}<11'b00111001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111001100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b00111001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00111001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111001111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b00111010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=11'b00111010001) && ({row_reg, col_reg}<11'b00111010100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111010100)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b00111010101)) color_data = 12'b101110101000;
		if(({row_reg, col_reg}==11'b00111010110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b00111011000) && ({row_reg, col_reg}<11'b00111011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111011100)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00111011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00111011110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00111011111)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=11'b00111100000) && ({row_reg, col_reg}<11'b00111100010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00111100010)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==11'b00111100011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00111100100)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b00111100101) && ({row_reg, col_reg}<11'b00111101000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111101000)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00111101001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00111101010)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00111101011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00111101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111101101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b00111101110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=11'b00111110000) && ({row_reg, col_reg}<11'b00111110011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111110011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b00111110100)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00111110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b00111110111)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==11'b00111111000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b00111111001)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b00111111010)) color_data = 12'b010100110010;

		if(({row_reg, col_reg}==11'b00111111011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01000000000) && ({row_reg, col_reg}<11'b01000000010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000000010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01000000011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01000000101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01000000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000000111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01000001000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01000001001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000001010)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}==11'b01000001011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000001100)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01000001101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01000001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000001111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01000010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=11'b01000010001) && ({row_reg, col_reg}<11'b01000010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000010110)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01000010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01000011000) && ({row_reg, col_reg}<11'b01000011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000011100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01000011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01000011110)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=11'b01000011111) && ({row_reg, col_reg}<11'b01000100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000100011)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==11'b01000100100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01000100101) && ({row_reg, col_reg}<11'b01000101000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000101000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01000101001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=11'b01000101010) && ({row_reg, col_reg}<11'b01000101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01000110000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01000110001) && ({row_reg, col_reg}<11'b01000110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000110100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01000110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01000110110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01000110111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000111000)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01000111001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01000111010)) color_data = 12'b011001000100;

		if(({row_reg, col_reg}==11'b01000111011)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01001000000) && ({row_reg, col_reg}<11'b01001000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001000101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01001000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001000111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01001001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b01001001001) && ({row_reg, col_reg}<11'b01001001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01001001101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01001001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001001111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01001010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01001010001)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b01001010010) && ({row_reg, col_reg}<11'b01001010100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001010100)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01001010101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001010110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01001010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01001011000) && ({row_reg, col_reg}<11'b01001011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001011100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01001011101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=11'b01001011110) && ({row_reg, col_reg}<11'b01001100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001100011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01001100100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01001100101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01001100110)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01001100111)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}==11'b01001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001101001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01001101010) && ({row_reg, col_reg}<11'b01001101101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001101101)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01001101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001101111)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01001110000)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==11'b01001110001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001110010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01001110011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001110100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01001110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01001110110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01001110111) && ({row_reg, col_reg}<11'b01001111001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01001111001)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==11'b01001111010)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==11'b01001111011)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01010000000) && ({row_reg, col_reg}<11'b01010000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010000101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01010000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010000111)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==11'b01010001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010001001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01010001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010001011)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==11'b01010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010001101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01010001110)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01010001111)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01010010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=11'b01010010001) && ({row_reg, col_reg}<11'b01010010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010010110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01010010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010011000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010011001)) color_data = 12'b110010101000;
		if(({row_reg, col_reg}>=11'b01010011010) && ({row_reg, col_reg}<11'b01010011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010011100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01010011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01010011110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01010011111) && ({row_reg, col_reg}<11'b01010100010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010100010)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01010100011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01010100100)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=11'b01010100101) && ({row_reg, col_reg}<11'b01010100111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010100111)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01010101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010101001)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}>=11'b01010101010) && ({row_reg, col_reg}<11'b01010101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010101100)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01010101101) && ({row_reg, col_reg}<11'b01010101111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010101111)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==11'b01010110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01010110001)) color_data = 12'b101110101000;
		if(({row_reg, col_reg}>=11'b01010110010) && ({row_reg, col_reg}<11'b01010110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010110100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01010110101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=11'b01010110110) && ({row_reg, col_reg}<11'b01010111001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01010111001)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01010111010)) color_data = 12'b011001010100;

		if(({row_reg, col_reg}==11'b01010111011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01011000000) && ({row_reg, col_reg}<11'b01011000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01011000101)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01011000110) && ({row_reg, col_reg}<11'b01011001000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01011001001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01011001010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011001011)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01011001100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b01011001101)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==11'b01011001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011001111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01011010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01011010001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011010010)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}>=11'b01011010011) && ({row_reg, col_reg}<11'b01011010101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011010101)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b01011010110)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==11'b01011010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01011011000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011011001)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}>=11'b01011011010) && ({row_reg, col_reg}<11'b01011011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011011100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01011011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01011011110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011011111)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b01011100000)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}>=11'b01011100001) && ({row_reg, col_reg}<11'b01011100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b01011100100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01011100101) && ({row_reg, col_reg}<11'b01011100111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011100111)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}==11'b01011101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01011101001)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01011101010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011101011)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01011101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011101101)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01011101110)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01011101111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01011110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01011110001)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01011110010) && ({row_reg, col_reg}<11'b01011110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011110100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01011110101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=11'b01011110110) && ({row_reg, col_reg}<11'b01011111000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01011111000)) color_data = 12'b110010111001;

		if(({row_reg, col_reg}>=11'b01011111001) && ({row_reg, col_reg}<11'b01100000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01100000101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01100000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100000111)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01100001000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01100001001)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==11'b01100001010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01100001011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01100001100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}>=11'b01100001101) && ({row_reg, col_reg}<11'b01100001111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100001111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01100010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01100010001)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}>=11'b01100010010) && ({row_reg, col_reg}<11'b01100010100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100010100)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b01100010101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100010110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01100010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01100011000) && ({row_reg, col_reg}<11'b01100011100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100011100)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==11'b01100011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b01100011110) && ({row_reg, col_reg}<11'b01100100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100100011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01100100100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01100100101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100100110)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01100100111)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}==11'b01100101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01100101001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01100101010) && ({row_reg, col_reg}<11'b01100101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100101110)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==11'b01100101111)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01100110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01100110001)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b01100110010) && ({row_reg, col_reg}<11'b01100110100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01100110100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01100110101)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}>=11'b01100110110) && ({row_reg, col_reg}<11'b01101000100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01101000101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01101000110)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01101000111)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101001000)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01101001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01101001010)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01101001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101001100)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==11'b01101001101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101001110)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01101001111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01101010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01101010001) && ({row_reg, col_reg}<11'b01101010110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101010110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01101010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01101011000) && ({row_reg, col_reg}<11'b01101011010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101011010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01101011011)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01101011100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01101011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01101011110) && ({row_reg, col_reg}<11'b01101100011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101100011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01101100100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01101100101) && ({row_reg, col_reg}<11'b01101101000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101101000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01101101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01101101010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101101011)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=11'b01101101100) && ({row_reg, col_reg}<11'b01101101110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101101110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101110000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b01101110001) && ({row_reg, col_reg}<11'b01101110011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01101110011)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==11'b01101110100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01101110101)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=11'b01101110110) && ({row_reg, col_reg}<11'b01110000000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110000000)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}==11'b01110000001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110000010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01110000011)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110000101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01110000110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110000111)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==11'b01110001000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110001001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01110001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01110001011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=11'b01110001100) && ({row_reg, col_reg}<11'b01110001110)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110001110)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01110001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01110010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110010001)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}>=11'b01110010010) && ({row_reg, col_reg}<11'b01110010101)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110010101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01110010110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01110010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110011000)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=11'b01110011001) && ({row_reg, col_reg}<11'b01110011011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110011011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01110011100)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01110011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01110011110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=11'b01110011111) && ({row_reg, col_reg}<11'b01110100010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110100010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01110100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=11'b01110100101) && ({row_reg, col_reg}<11'b01110101000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110101000)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==11'b01110101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01110101010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b01110101011)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01110101100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110101101)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=11'b01110101110) && ({row_reg, col_reg}<11'b01110110000)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=11'b01110110000) && ({row_reg, col_reg}<11'b01110110010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110110010)) color_data = 12'b110110101001;
		if(({row_reg, col_reg}==11'b01110110011)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110110100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01110110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01110110110)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=11'b01110110111) && ({row_reg, col_reg}<11'b01110111001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01110111001)) color_data = 12'b110110101001;

		if(({row_reg, col_reg}>=11'b01110111010) && ({row_reg, col_reg}<11'b01111000001)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111000001)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01111000010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01111000011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01111000100)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}>=11'b01111000101) && ({row_reg, col_reg}<11'b01111000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111000111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01111001000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111001001)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01111001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==11'b01111001011)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01111001100)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111001101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01111001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=11'b01111001111) && ({row_reg, col_reg}<11'b01111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111010010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01111010011)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==11'b01111010100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01111010101) && ({row_reg, col_reg}<11'b01111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111010111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111011000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01111011001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01111011010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01111011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01111011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111011101)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==11'b01111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111100001)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01111100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01111100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01111100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111100110)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01111100111) && ({row_reg, col_reg}<11'b01111101010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111101010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==11'b01111101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01111101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111101101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01111101110)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01111101111) && ({row_reg, col_reg}<11'b01111110010)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==11'b01111110010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==11'b01111110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b01111110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111110101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==11'b01111110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01111110111)) color_data = 12'b010101000011;





		if(({row_reg, col_reg}>=11'b01111111000) && ({row_reg, col_reg}<=11'b10011111011)) color_data = 12'b110010101001;
	end
endmodule